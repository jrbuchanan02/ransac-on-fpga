`timescale 1ns / 1ps

module derive_plane;
    // todo: place test here.
endmodule : derive_plane